module bubble(
    input clk,
    input rst,
    output b
);

endmodule