module wb(

);

endmodule